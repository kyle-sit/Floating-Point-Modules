/* File containing module code for a floating point multiplier
*/

//multiplier module
module multiplier_fp(
	input logic clk, start,
	input logic [31:0] A, B,
	output logic ready, busy,
	output logic [31:0] Y
);

endmodule